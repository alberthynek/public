LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Tape_Counter_TEST IS
	PORT(
			Clock, Reset, Increment, Decrement : IN STD_LOGIC;
			H1,H0,M1,M0,S1,S0 : OUT UNSIGNED (3 DOWNTO 0)
	);
END;

ARCHITECTURE behavioural OF Tape_Counter_TEST IS
	SIGNAL HH : UNSIGNED( 7 DOWNTO 0);
	SIGNAL MM : UNSIGNED( 7 DOWNTO 0);
	SIGNAL SS : UNSIGNED( 7 DOWNTO 0);
BEGIN
		PROCESS ( Clock )
		BEGIN 
			IF ( rising_edge (Clock)) THEN
				IF(Reset = '0')THEN
					HH <= "00";
					MM <= "00";
					SS <= "00";
				ELSIF ( Increment = '1') THEN
						IF (SS = "59") THEN
							SS <= "00";
							IF (MM = "59") THEN
								MM <= "00";
								IF (HH = "99") THEN
									HH <= "00";
								ELSE
									HH <= HH + 1;
								END IF;
							ELSE
								MM <= MM + 1;
							END IF;
						ELSE
							SS <= SS + 1;
						END IF;
				ELSIF ( Decrement = '1') THEN
						IF (SS = "00") THEN
							SS <= "59";
							IF (MM = "") THEN
								MM <= "59";
								IF (HH = "00") THEN
									HH <= "99";
								ELSE
									HH <= HH - 1;
								END IF;
							ELSE
								MM <= MM - 1;
							END IF;
						ELSE
							SS <= SS - 1;
						END IF;
				END IF;
			END IF;
		END PROCESS;
		
		H1 <= HH(7 DOWNTO 4);
		H0 <= HH(3 DOWNTO 0);
		M1 <= MM(7 DOWNTO 4);
		M0 <= MM(3 DOWNTO 0);
		S1 <= SS(7 DOWNTO 4);
		S0 <= SS(3 DOWNTO 0);
END;
						
						
							